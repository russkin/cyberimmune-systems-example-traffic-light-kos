component traffic_light.CReport

endpoints {
    report : traffic_light.IReport
}
